module osv

import time
import vlibuv
import vlibuv.uv

// FileInfo represents file metadata
pub struct FileInfo {
pub:
	path       string
	size       i64
	mode       u64
	uid        u32
	gid        u32
	atime      time.Time
	mtime      time.Time
	ctime      time.Time
	is_dir     bool
	is_file    bool
	is_link    bool
	is_fifo    bool
	is_socket  bool
	is_block   bool
	is_char    bool
}

// FileEvent represents a file system event
pub struct FileEvent {
pub:
	filename string
	events   int
	status   int
	is_rename bool
	is_change bool
}

// ============================================================================
// FILE OPERATIONS
// ============================================================================

// read_file reads the entire contents of a file
pub fn read_file(path string) ![]u8 {
	loop := vlibuv.Loop.default()

	// First, stat the file to get its size
	mut stat_req := uv.Uv_fs_t{}
	defer {
		uv.fs_req_cleanup(&stat_req)
	}

	// Synchronously stat the file
	uv.fs_stat(loop.get_c_loop(), &stat_req, path.str, fn (req &uv.Uv_fs_t) {})
	loop.run(uv.Mode.default)!

	stat_result := uv.fs_get_result(&stat_req)
	if stat_result < 0 {
		return error('failed to stat file: error code ${stat_result}')
	}

	// Get the file size from stat
	stat_buf := uv.fs_get_statbuf(&stat_req)
	if stat_buf == unsafe { nil } {
		return error('failed to get stat buffer')
	}

	file_size := 0 // TODO: Extract size from stat_buf when field is available

	// Open the file
	mut open_req := uv.Uv_fs_t{}
	defer {
		uv.fs_req_cleanup(&open_req)
	}

	uv.fs_open(loop.get_c_loop(), &open_req, path.str, 0, 0, fn (req &uv.Uv_fs_t) {})
	loop.run(uv.Mode.default)!

	fd := uv.fs_get_result(&open_req)
	if fd < 0 {
		return error('failed to open file: error code ${fd}')
	}

	// Allocate buffer for reading
	mut buffer := []u8{len: if file_size > 0 { file_size } else { 4096 }}

	// Read the file
	mut read_req := uv.Uv_fs_t{}
	defer {
		uv.fs_req_cleanup(&read_req)
	}

	// Create buf_t for reading - use data pointer of buffer
	buf := uv.buf_init(buffer.data, u32(buffer.len))

	uv.fs_read(loop.get_c_loop(), &read_req, fd, &buf, 1, 0, fn (req &uv.Uv_fs_t) {})
	loop.run(uv.Mode.default)!

	nread := uv.fs_get_result(&read_req)
	if nread < 0 {
		// Close file before returning error
		mut close_req := uv.Uv_fs_t{}
		defer {
			uv.fs_req_cleanup(&close_req)
		}
		uv.fs_close(loop.get_c_loop(), &close_req, fd, fn (req &uv.Uv_fs_t) {})
		loop.run(uv.Mode.default)!
		return error('failed to read file: error code ${nread}')
	}

	// Close the file
	mut close_req := uv.Uv_fs_t{}
	defer {
		uv.fs_req_cleanup(&close_req)
	}
	uv.fs_close(loop.get_c_loop(), &close_req, fd, fn (req &uv.Uv_fs_t) {})
	loop.run(uv.Mode.default)!

	return buffer[..nread]
}

// write_file writes data to a file, creating it if it doesn't exist
pub fn write_file(path string, data []u8) ! {
	loop := vlibuv.Loop.default()

	// Open file with create and write flags (0o644 = 420 in decimal)
	mut open_req := uv.Uv_fs_t{}
	defer {
		uv.fs_req_cleanup(&open_req)
	}

	flags := 0o666 | 0o1024 | 0o2000 // O_WRONLY | O_CREAT | O_TRUNC (approximate)
	uv.fs_open(loop.get_c_loop(), &open_req, path.str, flags, 0o644, fn (req &uv.Uv_fs_t) {})
	loop.run(uv.Mode.default)!

	fd := uv.fs_get_result(&open_req)
	if fd < 0 {
		return error('failed to open file for writing: error code ${fd}')
	}

	// Write data
	mut write_req := uv.Uv_fs_t{}
	defer {
		uv.fs_req_cleanup(&write_req)
	}

	buf := uv.buf_init(data.data, u32(data.len))

	uv.fs_write(loop.get_c_loop(), &write_req, fd, &buf, 1, 0, fn (req &uv.Uv_fs_t) {})
	loop.run(uv.Mode.default)!

	nwritten := uv.fs_get_result(&write_req)
	if nwritten < 0 {
		mut close_req := uv.Uv_fs_t{}
		defer {
			uv.fs_req_cleanup(&close_req)
		}
		uv.fs_close(loop.get_c_loop(), &close_req, fd, fn (req &uv.Uv_fs_t) {})
		loop.run(uv.Mode.default)!
		return error('failed to write file: error code ${nwritten}')
	}

	// Close the file
	mut close_req := uv.Uv_fs_t{}
	defer {
		uv.fs_req_cleanup(&close_req)
	}
	uv.fs_close(loop.get_c_loop(), &close_req, fd, fn (req &uv.Uv_fs_t) {})
	loop.run(uv.Mode.default)!
}

// append_file appends data to a file
pub fn append_file(path string, data []u8) ! {
	loop := vlibuv.Loop.default()

	// Open file with append and write flags
	mut open_req := uv.Uv_fs_t{}
	defer {
		uv.fs_req_cleanup(&open_req)
	}

	flags := 0o1 | 0o1024 | 0o10 // O_WRONLY | O_CREAT | O_APPEND (approximate)
	uv.fs_open(loop.get_c_loop(), &open_req, path.str, flags, 0o644, fn (req &uv.Uv_fs_t) {})
	loop.run(uv.Mode.default)!

	fd := uv.fs_get_result(&open_req)
	if fd < 0 {
		return error('failed to open file for appending: error code ${fd}')
	}

	// Write data
	mut write_req := uv.Uv_fs_t{}
	defer {
		uv.fs_req_cleanup(&write_req)
	}

	buf := uv.buf_init(data.data, u32(data.len))

	uv.fs_write(loop.get_c_loop(), &write_req, fd, &buf, 1, -1, fn (req &uv.Uv_fs_t) {})
	loop.run(uv.Mode.default)!

	nwritten := uv.fs_get_result(&write_req)
	if nwritten < 0 {
		mut close_req := uv.Uv_fs_t{}
		defer {
			uv.fs_req_cleanup(&close_req)
		}
		uv.fs_close(loop.get_c_loop(), &close_req, fd, fn (req &uv.Uv_fs_t) {})
		loop.run(uv.Mode.default)!
		return error('failed to append to file: error code ${nwritten}')
	}

	// Close the file
	mut close_req := uv.Uv_fs_t{}
	defer {
		uv.fs_req_cleanup(&close_req)
	}
	uv.fs_close(loop.get_c_loop(), &close_req, fd, fn (req &uv.Uv_fs_t) {})
	loop.run(uv.Mode.default)!
}

// remove_file deletes a file
pub fn remove_file(path string) ! {
	loop := vlibuv.Loop.default()

	mut req := uv.Uv_fs_t{}
	defer {
		uv.fs_req_cleanup(&req)
	}

	uv.fs_unlink(loop.get_c_loop(), &req, path.str, fn (req &uv.Uv_fs_t) {})
	loop.run(uv.Mode.default)!

	result := uv.fs_get_result(&req)
	if result < 0 {
		return error('failed to remove file: error code ${result}')
	}
}

// copy_file copies a file to a new location
pub fn copy_file(src string, dst string) ! {
	// Read the source file
	data := read_file(src)!
	// Write to destination
	write_file(dst, data)!
}

// rename_file renames or moves a file
pub fn rename_file(old_path string, new_path string) ! {
	loop := vlibuv.Loop.default()

	mut req := uv.Uv_fs_t{}
	defer {
		uv.fs_req_cleanup(&req)
	}

	uv.fs_rename(loop.get_c_loop(), &req, old_path.str, new_path.str, fn (req &uv.Uv_fs_t) {})
	loop.run(uv.Mode.default)!

	result := uv.fs_get_result(&req)
	if result < 0 {
		return error('failed to rename file: error code ${result}')
	}
}

// ============================================================================
// DIRECTORY OPERATIONS
// ============================================================================

// create_dir creates a directory
pub fn create_dir(path string, mode int) ! {
	// TODO: Implement using uv.fs_mkdir
}

// create_dir_all creates a directory and all parent directories
pub fn create_dir_all(path string, mode int) ! {
	// TODO: Implement creating parent directories
}

// remove_dir removes an empty directory
pub fn remove_dir(path string) ! {
	// TODO: Implement using uv.fs_rmdir
}

// DirEntry represents a directory entry
pub struct DirEntry {
pub:
	name    string
	is_file bool
	is_dir  bool
	is_link bool
}

// read_dir reads directory contents
pub fn read_dir(path string) ![]DirEntry {
	return []DirEntry{}
}

// ============================================================================
// FILE METADATA
// ============================================================================

// stat returns file information
pub fn stat(path string) !FileInfo {
	// TODO: Implement using uv.fs_stat
	return FileInfo{}
}

// lstat returns file information without following symlinks
pub fn lstat(path string) !FileInfo {
	// TODO: Implement using uv.fs_lstat
	return FileInfo{}
}

// exists checks if a file exists
pub fn exists(path string) bool {
	_ := stat(path) or { return false }
	return true
}

// is_file checks if path is a regular file
pub fn is_file(path string) bool {
	info := stat(path) or { return false }
	return info.is_file
}

// is_dir checks if path is a directory
pub fn is_dir(path string) bool {
	info := stat(path) or { return false }
	return info.is_dir
}

// is_link checks if path is a symlink
pub fn is_link(path string) bool {
	info := lstat(path) or { return false }
	return info.is_link
}

// ============================================================================
// SYMLINK & LINK OPERATIONS
// ============================================================================

// create_symlink creates a symbolic link
pub fn create_symlink(target string, linkpath string) ! {
	// TODO: Implement using uv.fs_symlink
}

// read_link reads the target of a symlink
pub fn read_link(path string) !string {
	// TODO: Implement using uv.fs_readlink
	return ''
}

// real_path returns the absolute path resolving symlinks
pub fn real_path(path string) !string {
	// TODO: Implement using uv.fs_realpath
	return ''
}

// create_hard_link creates a hard link
pub fn create_hard_link(target string, linkpath string) ! {
	// TODO: Implement using uv.fs_link
}

// ============================================================================
// FILE PERMISSIONS & OWNERSHIP
// ============================================================================

// chmod changes file permissions
pub fn chmod(path string, mode int) ! {
	// TODO: Implement using uv.fs_chmod
}

// fchmod changes permissions on an open file descriptor
pub fn fchmod(fd int, mode int) ! {
	// TODO: Implement using uv.fs_fchmod
}

// chown changes file owner and group
pub fn chown(path string, uid usize, gid usize) ! {
	// TODO: Implement using uv.fs_chown
}

// fchown changes ownership on an open file descriptor
pub fn fchown(fd int, uid usize, gid usize) ! {
	// TODO: Implement using uv.fs_fchown
}

// access checks file access permissions
pub fn access(path string, mode int) ! {
	// TODO: Implement using uv.fs_access
}

// ============================================================================
// FILE TIMES
// ============================================================================

// set_atime sets file access time
pub fn set_atime(path string, atime time.Time) ! {
	// TODO: Implement using uv.fs_utime
}

// set_mtime sets file modification time
pub fn set_mtime(path string, mtime time.Time) ! {
	// TODO: Implement using uv.fs_utime
}

// set_times sets both access and modification times
pub fn set_times(path string, atime time.Time, mtime time.Time) ! {
	// TODO: Implement using uv.fs_utime
}

// ============================================================================
// TEMPORARY FILES
// ============================================================================

// make_temp_dir creates a temporary directory
pub fn make_temp_dir(template string) !string {
	// TODO: Implement using uv.fs_mkdtemp
	return ''
}

// make_temp_file creates a temporary file
pub fn make_temp_file(template string) !(int, string) {
	// TODO: Implement using uv.fs_mkstemp
	return 0, ''
}

// ============================================================================
// FILE SYSTEM INFO
// ============================================================================

// StatFS holds file system statistics
pub struct StatFS {
pub:
	bsize   u64 // file system block size
	frsize  u64 // fragment size
	blocks  u64 // size of fs in frsize units
	bfree   u64 // # free blocks
	bavail  u64 // # free blocks for non-root
	files   u64 // # inodes
	ffree   u64 // # free inodes
	favail  u64 // # free inodes for non-root
	flag    u64 // mount flags
	namemax u64 // maximum filename length
}

// stat_fs returns file system statistics
pub fn stat_fs(path string) !StatFS {
	// TODO: Implement using uv.fs_statfs
	return StatFS{}
}

// ============================================================================
// FILE WATCHING
// ============================================================================

pub struct FileWatcher {
mut:
	handle   &uv.Uv_fs_event_t
	path     string
	callback ?fn(event FileEvent) = unsafe { nil }
	running  bool
}

// watch_file watches a file for changes
pub fn watch_file(path string, callback fn(event FileEvent)) !FileWatcher {
	return FileWatcher{
		handle: &uv.Uv_fs_event_t{}
		path: path
		callback: callback
		running: false
	}
}

// stop stops watching the file
pub fn (mut w FileWatcher) stop() ! {
	// TODO: Implement proper file watcher stop
	w.running = false
}
