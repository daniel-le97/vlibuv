module vlibuv

pub type Buf = C.uv_buf_t
