module vlibuv

// pub struct Work {
// 	Req // pub mut:
// 	// 	l_data voidptr = unsafe { nil }
// }

// pub fn new_work() Work {
// 	work := &C.uv_work_t(unsafe { nil })
// 	return Work{Req{work, unsafe { nil }}}
// }

// pub fn new_worker() &C.uv_work_t {
// 	work := &C.uv_work_t{}
// 	// work := &C.uv_work_t(unsafe { nil })
// 	return work
// }

// pub fn (w Work) to_work() &C.uv_work_t {
// 	unsafe {
// 		return &C.uv_work_t(w.req)
// 	}
// }
