module vuv
