module vlibuv
