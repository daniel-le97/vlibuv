module vlibuv

struct Work {
	Req

}





